					----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:27:38 02/16/2011 
-- Design Name: 
-- Module Name:    input_ctr - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity x4_input_ctr is
    Port ( clk : 					in  STD_LOGIC;
           init : 				in  STD_LOGIC;
           init_ev : 			in  STD_LOGIC;
			  wr_fifo_vme : 			in  STD_LOGIC;									--write enable of FIF
			  vme_input_fifo : 	in  STD_LOGIC_VECTOR (19 downto 0);		--hit in input of FIFO  
			  new_hit : 			in  STD_LOGIC;									--register enable of hit from P3
           lay_in :	 			in  STD_LOGIC_VECTOR (17 downto 0);		--hit in input from P3  
			  wr_hit_lamb :		in  STD_LOGIC;									--register nable of hit to lamb
			  hitmask : 			in  STD_LOGIC_VECTOR (17 downto 0);		--mask of hit		
			  tmode : 				in  STD_LOGIC;									--test mode (read each event from FIFO)
           edro_mode : 			in  STD_LOGIC;									--psuh out the hit from P3 connector
           start_rd_fifo : 	in  STD_LOGIC;									--start the read of FIFO when it's finish to write 
			  state  : 				in  STD_LOGIC_VECTOR (2 downto 0);		--current state of FSM
			  hit_loop  : 			in  STD_LOGIC;
			  
			  vmedata : 			in  STD_LOGIC_VECTOR (31 downto 0);
			  wr_nloop : 			in  STD_LOGIC;
			  			  
			  rd_fifo : 		out  STD_LOGIC;								--read fifo of hit
			  hee_reg : 		buffer  STD_LOGIC; 								--end event register
			  tag_ee_word :  	out  STD_LOGIC_VECTOR (15 downto 0);	--word of end event
        A_HIT : 			out  STD_LOGIC_VECTOR (17 downto 0);
			  enA_wr :			out  STD_LOGIC;			
			  HIT_lay : 		out  STD_LOGIC_VECTOR (17 downto 0);		--copy of hit in input (AMBSlim2)
			  push_hit : 		out  STD_LOGIC;									--data stobe of hit copy		  
			  data_ispy : 			buffer STD_LOGIC_VECTOR (20 downto 0);		--data storage in the ispy buffer
			  push_data_ispy : 	out STD_LOGIC									--data stobe of hit in the ispy buffer		  
			  
			  );
end x4_input_ctr;

architecture Behavioral of x4_input_ctr is
		
		--istanziate the fifo that storage the input write from VME
		component hit_fifo_vme is 
							port (clk: IN std_logic;
									rst: IN std_logic;
									din: IN std_logic_VECTOR(17 downto 0);
									wr_en: IN std_logic;
									rd_en: IN std_logic;
									dout: OUT std_logic_VECTOR(17 downto 0);
									full: OUT std_logic;
									empty: OUT std_logic
									);
		end component hit_fifo_vme;
		
		--input hit register
		signal lay_reg : STD_LOGIC_VECTOR (17 downto 0);
		
		--signal of fifo
		signal empty_fifo : STD_LOGIC;
		signal rd_fifo_edro_mode : STD_LOGIC;
		signal rd_fifo_tmode : STD_LOGIC;
		signal rd_en_reg : STD_LOGIC;
		
		--end event in out of FIFO
		signal ee_out_fifo : STD_LOGIC;
		
		--data in input at the register before the output
		signal data : STD_LOGIC_VECTOR (17 downto 0);
		
		--signal out from FIFO
		signal vme_out_fifo : STD_LOGIC_VECTOR (17 downto 0);
		
		signal vme_reg : STD_LOGIC_VECTOR (17 downto 0);
		
		--this signal is an input generated by FSM
		signal rd_fifo_int : STD_LOGIC;
		signal rd_fifo_d1 : STD_LOGIC;
		
		--this signal is usefull when the FSM is in the 3 state
		signal state3 : STD_LOGIC;
		signal new_event_d1 : STD_LOGIC;
		
		--signal of FIFO
		signal data_input_fifo : STD_LOGIC_VECTOR (17 downto 0);
		signal wr_fifo_loop : STD_LOGIC;
		signal wr_fifo : STD_LOGIC;
		
		--data ispy
		signal push_ispy : STD_LOGIC;
		
		--signal to register the counter of number the loop of fifo
		signal wr_nloop_d1 : STD_LOGIC;
		signal wr_nloop_d2 : STD_LOGIC;
		signal wr_nloop_d3 : STD_LOGIC;
		signal wr_nloop_pulse : STD_LOGIC;
		signal wr_pulse_comp : STD_LOGIC;
		
		--signal to enable the counter
		signal en_counter : STD_LOGIC;
		signal en_counter_d1 : STD_LOGIC;
		signal en_counter_d2 : STD_LOGIC;
		
		
		signal mask_loop : STD_LOGIC;
		signal event_zero : STD_LOGIC;
		signal zero_loop : STD_LOGIC;
		
		--value of the loop number of the FIFO
		signal counter_nloop : STD_LOGIC_VECTOR (31 downto 0);
		
		
		
begin
		
		--signal to create the loop of the FIFO
		data_input_fifo <= vme_out_fifo when hit_loop = '1' else vme_input_fifo(17 downto 0);
		
		wr_fifo <= wr_fifo_loop when hit_loop = '1' else wr_fifo_vme;
		
		wr_fifo_loop <= rd_fifo_d1 and mask_loop;
		
				--control if the counter is zero to determinate a infinite loop
		comparator_proc: process(clk, init)
		begin
			if(init = '1') then
				zero_loop <= '0';
			elsif(clk'event and clk = '1') then
				if(wr_pulse_comp = '1' and counter_nloop = "00000000000000000000000000000000") then
					zero_loop <= '1';
				end if;
			end if;
		end process;
		
		wr_pulse_comp <= (not wr_nloop_d3) and wr_nloop_d2;
		--define the process to create a pulse to storage the value of the counter
		--in the register adressed by VME
		wr_nloop_proc : process(clk, init)
		begin
			if(init = '1') then
				wr_nloop_d1 <= '0';
				wr_nloop_d2 <= '0';
			elsif(clk'event and clk = '1') then
				wr_nloop_d1 <= wr_nloop;
				wr_nloop_d2 <= wr_nloop_d1;
				wr_nloop_d3 <= wr_nloop_d2;
			end if;
		end process;
		
		wr_nloop_pulse <= (not wr_nloop_d2) and wr_nloop_d1;
		
		--comparator of event number zero
		event_zero <= '1' when vme_out_fifo(15 downto 0) = "0000000000000000" else '0';
		
		--enable the counter if the value of counter id not zero; if there is the 
		--loop mode; if there is the event zero and the mask is enable
		--en_counter <= (not zero_loop) and event_zero and hit_loop and mask_loop and rd_fifo_d1;
		en_counter <= (not zero_loop) and event_zero and hit_loop and wr_fifo_loop;
		
		en_counter_proc : process(clk, init)
		begin
			if(init = '1') then
				en_counter_d1 <= '0';
				en_counter_d2 <= '0';
			elsif(clk'event and clk = '1') then
					en_counter_d1 <= en_counter;
					en_counter_d2 <= en_counter_d1;
			end if;
		end process;
				
	
		--register the value of the counter and count the nummber of cycle of the FIFO
		couter_process: process(clk, init)
		begin
			if(init = '1') then
				mask_loop <= '1';					--precharge the mask_loop at 1 
				counter_nloop <= "00000000000000000000000000000000";
			elsif(clk'event and clk = '1') then
				if(wr_nloop_pulse = '1') then		--storage the value of the counter
					counter_nloop <= vmedata;
				elsif(en_counter_d2 = '1') then
					counter_nloop <= counter_nloop - 1;
				elsif(counter_nloop = "00000000000000000000000000000000" and en_counter_d1 = '1') then
					mask_loop <= '0';
				end if;
			end if;
		end process;

		--the FIFO that storage the hit write from VME 
		--we can take all time to storage the hit 
		fifo: hit_fifo_vme port map(	clk => clk,
												rst => init,
												din => data_input_fifo,
												wr_en => wr_fifo,
												rd_en => rd_fifo_int,
												dout => vme_out_fifo,
												--full =>
												empty => empty_fifo
											);
		
		--control the bit of end event in out of FIFO
		ee_out_fifo <= vme_out_fifo(16);
		
		--logic to read FIFO when it's not empty and it's set the register to
		--give the start of read the fifo
		--when there is the word of end event in output of FIFO we can stop the read
		--of FIFO and restart when the FSM is in the state 3 (the cysle of event is finished)
		--and there is a new event
		rd_fifo_tmode <= start_rd_fifo and (not empty_fifo) and (new_event_d1 or not(ee_out_fifo));
		
		--consider the signal of state 3 to restart the read of FIFO
		state3 <= '1' when state="111" else '0';
		
		process(clk, init)
		begin
			if(init = '1') then
				new_event_d1 <= '0';
			elsif(clk'event and clk='1') then
				new_event_d1 <= state3;
			end if;
		end process;
		
		--select the mode of run. If it's in EDRO mode we can push out the hit 
		-- and the control is the signal empty; when i's in test mode the read
		--of FIFO is control by the logic 
		rd_fifo_int <= rd_fifo_edro_mode when edro_mode = '1' else rd_fifo_tmode;
		
		--signal to enable the register
		process(clk)
		begin
			if(clk'event and clk='1') then
				rd_en_reg <= rd_fifo_int;
			end if;
		end process;
		
		--assign the signal of read fifo in output
		rd_fifo <= rd_fifo_int;
			
		--insert the register for the data in output of FIFO
		process (clk, init, init_ev)
		begin
			if (init = '1' or init_ev ='1') then
				vme_reg <= (others => '0');
			elsif (clk'event and clk = '1') then
				if (rd_en_reg = '1') then
					vme_reg <= vme_out_fifo;
				end if;
			end if;
		end process;
		
		--register the hit in input for normal mode
		process (clk, init, init_ev)
		begin
			if (init = '1' or init_ev = '1') then
				lay_reg <= (others => '0');
			elsif (clk'event and clk = '1') then
				if (new_hit = '1') then
					lay_reg <= lay_in(17 downto 0);
				end if;
			end if;
		end process;
		
		
		--mux to select the mode of run
		data <= lay_reg(17 downto 0) when tmode = '0' else vme_reg(17 downto 0);
		
		--signal to write the hit in ispy
		data_ispy <= ("000" & data);
		
		push_ispy <= new_hit when tmode='0' else rd_en_reg;
		
		process(clk)
		begin
			if(clk'event and clk='1')then
				push_data_ispy <= push_ispy;
			end if;
		end process;
		
		--define the tag of each event
		process (clk, init)
		begin
			if (init = '1') then
				tag_ee_word <= (others => '0');
			elsif(clk'event and clk = '1') then
				if(data(16) = '1') then
					tag_ee_word <= data(15 downto 0);
				end if;
			end if;
		end process;
		
		--assign the end event 
		hee_reg <= data(16);

		--register the hit before the output of chip
		process (clk, init_ev)
		begin
			if (init_ev = '1') then
				A_HIT <= (others => '0');
			elsif (clk'event and clk = '1') then
				if(wr_hit_lamb = '1') then
					A_HIT <= (data or hitmask);
				end if;
			end if;
		end process;
		
		--data strobe for hit to lamb
		process(clk, init_ev)
		begin
			if(init_ev = '1') then
-- Guido - Nov 22
--				enA_wr <= '1';
--				enB_wr <= '1';
--				enC_wr <= '1';
--				enD_wr <= '1';
				enA_wr <= '0';
			elsif(clk'event and clk = '1') then
				enA_wr <= wr_hit_lamb;
			end if;
		end process;
		
		
		--******************************************************************
		--EDRO MODE
		--read FIFO in EDRO mode
		rd_fifo_edro_mode <= start_rd_fifo and (not empty_fifo);
		
		--register the hit before send out from P3
		--se serve l'abilitazione possiamo mettere il rd_fifo ri
		process (clk, init)
		begin
			if (init = '1') then
				HIT_lay <= (others => '0');
			elsif (clk'event and clk = '1') then
				HIT_lay <= vme_out_fifo;
			end if;
		end process;
		
		--data stobe of hit in out
		process (clk, init)
		begin
			if (init = '1') then
				rd_fifo_d1 <= '0';
				push_hit <= '0';
			elsif(clk'event and clk = '1') then
				rd_fifo_d1 <= rd_fifo_int;
				push_hit <= rd_fifo_d1;
			end if;
		end process;

	
end Behavioral;

